module and_gate(
    input a,
    input b,
    output z
    );
  assign z = ~(a | b);

endmodule
